** Profile: "SCHEMATIC1-dioda"  [ c:\users\coste\onedrive\desktop\cad\lab5-pspicefiles\proiect cad-PSpiceFiles\SCHEMATIC1\dioda.sim ] 

** Creating circuit file "dioda.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Users\coste\OneDrive\Desktop\an2\sem2\workspace_orcad\cdssetup\OrCAD_PSpice\23.1.0\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 1000ns 0 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
