** Profile: "SCHEMATIC1-tranzistor"  [ c:\users\coste\onedrive\desktop\cad\lab5-pspicefiles\proiect cad-PSpiceFiles\SCHEMATIC1\tranzistor.sim ] 

** Creating circuit file "tranzistor.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Users\coste\OneDrive\Desktop\an2\sem2\workspace_orcad\cdssetup\OrCAD_PSpice\23.1.0\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.DC LIN V_V4 -10 10 0.01 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
